----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:09:26 11/11/2021 
-- Design Name: 
-- Module Name:    top - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity top is
    Port ( M1 : in  STD_LOGIC;
           M2 : in  STD_LOGIC;
           M3 : in  STD_LOGIC;
           M4 : in  STD_LOGIC;
           N1 : in  STD_LOGIC;
           N2 : in  STD_LOGIC;
           N3 : in  STD_LOGIC;
           N4 : in  STD_LOGIC;
           START : in  STD_LOGIC;
           R1 : out  STD_LOGIC;
           R2 : out  STD_LOGIC;
           R3 : out  STD_LOGIC;
           R4 : out  STD_LOGIC;
           R5 : out  STD_LOGIC;
           R6 : out  STD_LOGIC;
           R7 : out  STD_LOGIC;
           R8 : out  STD_LOGIC;
           DONE : out  STD_LOGIC);
end top;

architecture Behavioral of top is

begin


end Behavioral;

